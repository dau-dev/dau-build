`timescale 1ns/1ns

module priorityencoder #(parameter SIZE = 5) (
	input logic [2**SIZE-1:0] inp_i,
	output logic [SIZE-1:0] out_o,
	output logic valid_o
);


always_comb begin
	casez (inp_i)
		32'b0000_0000_0000_0000_0000_0000_0000_0001: out_o=5'd0;
		32'b0000_0000_0000_0000_0000_0000_0000_001?: out_o=5'd1;
		32'b0000_0000_0000_0000_0000_0000_0000_01??: out_o=5'd2;
		32'b0000_0000_0000_0000_0000_0000_0000_1???: out_o=5'd3;
		32'b0000_0000_0000_0000_0000_0000_0001_????: out_o=5'd4;
		32'b0000_0000_0000_0000_0000_0000_001?_????: out_o=5'd5;
		32'b0000_0000_0000_0000_0000_0000_01??_????: out_o=5'd6;
		32'b0000_0000_0000_0000_0000_0000_1???_????: out_o=5'd7;
		32'b0000_0000_0000_0000_0000_0001_????_????: out_o=5'd8;
		32'b0000_0000_0000_0000_0000_001?_????_????: out_o=5'd9;
		32'b0000_0000_0000_0000_0000_01??_????_????: out_o=5'd10;
		32'b0000_0000_0000_0000_0000_1???_????_????: out_o=5'd11;
		32'b0000_0000_0000_0000_0001_????_????_????: out_o=5'd12;
		32'b0000_0000_0000_0000_001?_????_????_????: out_o=5'd13;
		32'b0000_0000_0000_0000_01??_????_????_????: out_o=5'd14;
		32'b0000_0000_0000_0000_1???_????_????_????: out_o=5'd15;
		32'b0000_0000_0000_0001_????_????_????_????: out_o=5'd16;
		32'b0000_0000_0000_001?_????_????_????_????: out_o=5'd17;
		32'b0000_0000_0000_01??_????_????_????_????: out_o=5'd18;
		32'b0000_0000_0000_1???_????_????_????_????: out_o=5'd19;
		32'b0000_0000_0001_????_????_????_????_????: out_o=5'd20;
		32'b0000_0000_001?_????_????_????_????_????: out_o=5'd21;
		32'b0000_0000_01??_????_????_????_????_????: out_o=5'd22;
		32'b0000_0000_1???_????_????_????_????_????: out_o=5'd23;
		32'b0000_0001_????_????_????_????_????_????: out_o=5'd24;
		32'b0000_001?_????_????_????_????_????_????: out_o=5'd25;
		32'b0000_01??_????_????_????_????_????_????: out_o=5'd26;
		32'b0000_1???_????_????_????_????_????_????: out_o=5'd27;
		32'b0001_????_????_????_????_????_????_????: out_o=5'd28;
		32'b001?_????_????_????_????_????_????_????: out_o=5'd29;
		32'b01??_????_????_????_????_????_????_????: out_o=5'd30;
		32'b1???_????_????_????_????_????_????_????: out_o=5'd31;
	endcase

	if (inp_i == 32'd0) begin
		valid_o = 1'b0;
	end

	else begin
		valid_o = 1'b1;
	end
end

endmodule
